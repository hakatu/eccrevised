  // polynomial: x^8 + x^2 + x^1 + 1
  // data width: 256
  // convention: the first serial bit is D[255]

module crc8_256
    (
     idat,
     icrc,
     ocrc
     );
input [255:0] idat;
input [7:0]   icrc;
output [7:0]  ocrc;

assign        ocrc[0] = idat[254]^idat[246]^idat[245]^idat[243]^idat[242]^idat[240]^idat[239]^idat[238]^idat[237]^idat[234]^idat[233]^idat[232]^idat[231]^idat[230]^idat[229]^idat[227]^idat[224]^idat[221]^idat[220]^idat[219]^idat[217]^idat[215]^idat[214]^idat[213]^idat[212]^idat[211]^idat[207]^idat[204]^idat[202]^idat[201]^idat[196]^idat[195]^idat[194]^idat[193]^idat[191]^idat[190]^idat[187]^idat[183]^idat[181]^idat[180]^idat[179]^idat[177]^idat[176]^idat[175]^idat[172]^idat[170]^idat[167]^idat[166]^idat[162]^idat[161]^idat[158]^idat[157]^idat[155]^idat[150]^idat[148]^idat[146]^idat[145]^idat[143]^idat[141]^idat[139]^idat[135]^idat[134]^idat[133]^idat[127]^idat[119]^idat[118]^idat[116]^idat[115]^idat[113]^idat[112]^idat[111]^idat[110]^idat[107]^idat[106]^idat[105]^idat[104]^idat[103]^idat[102]^idat[100]^idat[97]^idat[94]^idat[93]^idat[92]^idat[90]^idat[88]^idat[87]^idat[86]^idat[85]^idat[84]^idat[80]^idat[77]^idat[75]^idat[74]^idat[69]^idat[68]^idat[67]^idat[66]^idat[64]^idat[63]^idat[60]^idat[56]^idat[54]^idat[53]^idat[52]^idat[50]^idat[49]^idat[48]^idat[45]^idat[43]^idat[40]^idat[39]^idat[35]^idat[34]^idat[31]^idat[30]^idat[28]^idat[23]^idat[21]^idat[19]^idat[18]^idat[16]^idat[14]^idat[12]^idat[8]^idat[7]^idat[6]^idat[0]^icrc[6];
assign        ocrc[1] = idat[255]^idat[254]^idat[247]^idat[245]^idat[244]^idat[242]^idat[241]^idat[237]^idat[235]^idat[229]^idat[228]^idat[227]^idat[225]^idat[224]^idat[222]^idat[219]^idat[218]^idat[217]^idat[216]^idat[211]^idat[208]^idat[207]^idat[205]^idat[204]^idat[203]^idat[201]^idat[197]^idat[193]^idat[192]^idat[190]^idat[188]^idat[187]^idat[184]^idat[183]^idat[182]^idat[179]^idat[178]^idat[175]^idat[173]^idat[172]^idat[171]^idat[170]^idat[168]^idat[166]^idat[163]^idat[161]^idat[159]^idat[157]^idat[156]^idat[155]^idat[151]^idat[150]^idat[149]^idat[148]^idat[147]^idat[145]^idat[144]^idat[143]^idat[142]^idat[141]^idat[140]^idat[139]^idat[136]^idat[133]^idat[128]^idat[127]^idat[120]^idat[118]^idat[117]^idat[115]^idat[114]^idat[110]^idat[108]^idat[102]^idat[101]^idat[100]^idat[98]^idat[97]^idat[95]^idat[92]^idat[91]^idat[90]^idat[89]^idat[84]^idat[81]^idat[80]^idat[78]^idat[77]^idat[76]^idat[74]^idat[70]^idat[66]^idat[65]^idat[63]^idat[61]^idat[60]^idat[57]^idat[56]^idat[55]^idat[52]^idat[51]^idat[48]^idat[46]^idat[45]^idat[44]^idat[43]^idat[41]^idat[39]^idat[36]^idat[34]^idat[32]^idat[30]^idat[29]^idat[28]^idat[24]^idat[23]^idat[22]^idat[21]^idat[20]^idat[18]^idat[17]^idat[16]^idat[15]^idat[14]^idat[13]^idat[12]^idat[9]^idat[6]^idat[1]^idat[0]^icrc[6]^icrc[7];
assign        ocrc[2] = idat[255]^idat[254]^idat[248]^idat[240]^idat[239]^idat[237]^idat[236]^idat[234]^idat[233]^idat[232]^idat[231]^idat[228]^idat[227]^idat[226]^idat[225]^idat[224]^idat[223]^idat[221]^idat[218]^idat[215]^idat[214]^idat[213]^idat[211]^idat[209]^idat[208]^idat[207]^idat[206]^idat[205]^idat[201]^idat[198]^idat[196]^idat[195]^idat[190]^idat[189]^idat[188]^idat[187]^idat[185]^idat[184]^idat[181]^idat[177]^idat[175]^idat[174]^idat[173]^idat[171]^idat[170]^idat[169]^idat[166]^idat[164]^idat[161]^idat[160]^idat[156]^idat[155]^idat[152]^idat[151]^idat[149]^idat[144]^idat[142]^idat[140]^idat[139]^idat[137]^idat[135]^idat[133]^idat[129]^idat[128]^idat[127]^idat[121]^idat[113]^idat[112]^idat[110]^idat[109]^idat[107]^idat[106]^idat[105]^idat[104]^idat[101]^idat[100]^idat[99]^idat[98]^idat[97]^idat[96]^idat[94]^idat[91]^idat[88]^idat[87]^idat[86]^idat[84]^idat[82]^idat[81]^idat[80]^idat[79]^idat[78]^idat[74]^idat[71]^idat[69]^idat[68]^idat[63]^idat[62]^idat[61]^idat[60]^idat[58]^idat[57]^idat[54]^idat[50]^idat[48]^idat[47]^idat[46]^idat[44]^idat[43]^idat[42]^idat[39]^idat[37]^idat[34]^idat[33]^idat[29]^idat[28]^idat[25]^idat[24]^idat[22]^idat[17]^idat[15]^idat[13]^idat[12]^idat[10]^idat[8]^idat[6]^idat[2]^idat[1]^idat[0]^icrc[0]^icrc[6]^icrc[7];
assign        ocrc[3] = idat[255]^idat[249]^idat[241]^idat[240]^idat[238]^idat[237]^idat[235]^idat[234]^idat[233]^idat[232]^idat[229]^idat[228]^idat[227]^idat[226]^idat[225]^idat[224]^idat[222]^idat[219]^idat[216]^idat[215]^idat[214]^idat[212]^idat[210]^idat[209]^idat[208]^idat[207]^idat[206]^idat[202]^idat[199]^idat[197]^idat[196]^idat[191]^idat[190]^idat[189]^idat[188]^idat[186]^idat[185]^idat[182]^idat[178]^idat[176]^idat[175]^idat[174]^idat[172]^idat[171]^idat[170]^idat[167]^idat[165]^idat[162]^idat[161]^idat[157]^idat[156]^idat[153]^idat[152]^idat[150]^idat[145]^idat[143]^idat[141]^idat[140]^idat[138]^idat[136]^idat[134]^idat[130]^idat[129]^idat[128]^idat[122]^idat[114]^idat[113]^idat[111]^idat[110]^idat[108]^idat[107]^idat[106]^idat[105]^idat[102]^idat[101]^idat[100]^idat[99]^idat[98]^idat[97]^idat[95]^idat[92]^idat[89]^idat[88]^idat[87]^idat[85]^idat[83]^idat[82]^idat[81]^idat[80]^idat[79]^idat[75]^idat[72]^idat[70]^idat[69]^idat[64]^idat[63]^idat[62]^idat[61]^idat[59]^idat[58]^idat[55]^idat[51]^idat[49]^idat[48]^idat[47]^idat[45]^idat[44]^idat[43]^idat[40]^idat[38]^idat[35]^idat[34]^idat[30]^idat[29]^idat[26]^idat[25]^idat[23]^idat[18]^idat[16]^idat[14]^idat[13]^idat[11]^idat[9]^idat[7]^idat[3]^idat[2]^idat[1]^icrc[1]^icrc[7];
assign        ocrc[4] = idat[250]^idat[242]^idat[241]^idat[239]^idat[238]^idat[236]^idat[235]^idat[234]^idat[233]^idat[230]^idat[229]^idat[228]^idat[227]^idat[226]^idat[225]^idat[223]^idat[220]^idat[217]^idat[216]^idat[215]^idat[213]^idat[211]^idat[210]^idat[209]^idat[208]^idat[207]^idat[203]^idat[200]^idat[198]^idat[197]^idat[192]^idat[191]^idat[190]^idat[189]^idat[187]^idat[186]^idat[183]^idat[179]^idat[177]^idat[176]^idat[175]^idat[173]^idat[172]^idat[171]^idat[168]^idat[166]^idat[163]^idat[162]^idat[158]^idat[157]^idat[154]^idat[153]^idat[151]^idat[146]^idat[144]^idat[142]^idat[141]^idat[139]^idat[137]^idat[135]^idat[131]^idat[130]^idat[129]^idat[123]^idat[115]^idat[114]^idat[112]^idat[111]^idat[109]^idat[108]^idat[107]^idat[106]^idat[103]^idat[102]^idat[101]^idat[100]^idat[99]^idat[98]^idat[96]^idat[93]^idat[90]^idat[89]^idat[88]^idat[86]^idat[84]^idat[83]^idat[82]^idat[81]^idat[80]^idat[76]^idat[73]^idat[71]^idat[70]^idat[65]^idat[64]^idat[63]^idat[62]^idat[60]^idat[59]^idat[56]^idat[52]^idat[50]^idat[49]^idat[48]^idat[46]^idat[45]^idat[44]^idat[41]^idat[39]^idat[36]^idat[35]^idat[31]^idat[30]^idat[27]^idat[26]^idat[24]^idat[19]^idat[17]^idat[15]^idat[14]^idat[12]^idat[10]^idat[8]^idat[4]^idat[3]^idat[2]^icrc[2];
assign        ocrc[5] = idat[251]^idat[243]^idat[242]^idat[240]^idat[239]^idat[237]^idat[236]^idat[235]^idat[234]^idat[231]^idat[230]^idat[229]^idat[228]^idat[227]^idat[226]^idat[224]^idat[221]^idat[218]^idat[217]^idat[216]^idat[214]^idat[212]^idat[211]^idat[210]^idat[209]^idat[208]^idat[204]^idat[201]^idat[199]^idat[198]^idat[193]^idat[192]^idat[191]^idat[190]^idat[188]^idat[187]^idat[184]^idat[180]^idat[178]^idat[177]^idat[176]^idat[174]^idat[173]^idat[172]^idat[169]^idat[167]^idat[164]^idat[163]^idat[159]^idat[158]^idat[155]^idat[154]^idat[152]^idat[147]^idat[145]^idat[143]^idat[142]^idat[140]^idat[138]^idat[136]^idat[132]^idat[131]^idat[130]^idat[124]^idat[116]^idat[115]^idat[113]^idat[112]^idat[110]^idat[109]^idat[108]^idat[107]^idat[104]^idat[103]^idat[102]^idat[101]^idat[100]^idat[99]^idat[97]^idat[94]^idat[91]^idat[90]^idat[89]^idat[87]^idat[85]^idat[84]^idat[83]^idat[82]^idat[81]^idat[77]^idat[74]^idat[72]^idat[71]^idat[66]^idat[65]^idat[64]^idat[63]^idat[61]^idat[60]^idat[57]^idat[53]^idat[51]^idat[50]^idat[49]^idat[47]^idat[46]^idat[45]^idat[42]^idat[40]^idat[37]^idat[36]^idat[32]^idat[31]^idat[28]^idat[27]^idat[25]^idat[20]^idat[18]^idat[16]^idat[15]^idat[13]^idat[11]^idat[9]^idat[5]^idat[4]^idat[3]^icrc[3];
assign        ocrc[6] = idat[252]^idat[244]^idat[243]^idat[241]^idat[240]^idat[238]^idat[237]^idat[236]^idat[235]^idat[232]^idat[231]^idat[230]^idat[229]^idat[228]^idat[227]^idat[225]^idat[222]^idat[219]^idat[218]^idat[217]^idat[215]^idat[213]^idat[212]^idat[211]^idat[210]^idat[209]^idat[205]^idat[202]^idat[200]^idat[199]^idat[194]^idat[193]^idat[192]^idat[191]^idat[189]^idat[188]^idat[185]^idat[181]^idat[179]^idat[178]^idat[177]^idat[175]^idat[174]^idat[173]^idat[170]^idat[168]^idat[165]^idat[164]^idat[160]^idat[159]^idat[156]^idat[155]^idat[153]^idat[148]^idat[146]^idat[144]^idat[143]^idat[141]^idat[139]^idat[137]^idat[133]^idat[132]^idat[131]^idat[125]^idat[117]^idat[116]^idat[114]^idat[113]^idat[111]^idat[110]^idat[109]^idat[108]^idat[105]^idat[104]^idat[103]^idat[102]^idat[101]^idat[100]^idat[98]^idat[95]^idat[92]^idat[91]^idat[90]^idat[88]^idat[86]^idat[85]^idat[84]^idat[83]^idat[82]^idat[78]^idat[75]^idat[73]^idat[72]^idat[67]^idat[66]^idat[65]^idat[64]^idat[62]^idat[61]^idat[58]^idat[54]^idat[52]^idat[51]^idat[50]^idat[48]^idat[47]^idat[46]^idat[43]^idat[41]^idat[38]^idat[37]^idat[33]^idat[32]^idat[29]^idat[28]^idat[26]^idat[21]^idat[19]^idat[17]^idat[16]^idat[14]^idat[12]^idat[10]^idat[6]^idat[5]^idat[4]^icrc[4];
assign        ocrc[7] = idat[253]^idat[245]^idat[244]^idat[242]^idat[241]^idat[239]^idat[238]^idat[237]^idat[236]^idat[233]^idat[232]^idat[231]^idat[230]^idat[229]^idat[228]^idat[226]^idat[223]^idat[220]^idat[219]^idat[218]^idat[216]^idat[214]^idat[213]^idat[212]^idat[211]^idat[210]^idat[206]^idat[203]^idat[201]^idat[200]^idat[195]^idat[194]^idat[193]^idat[192]^idat[190]^idat[189]^idat[186]^idat[182]^idat[180]^idat[179]^idat[178]^idat[176]^idat[175]^idat[174]^idat[171]^idat[169]^idat[166]^idat[165]^idat[161]^idat[160]^idat[157]^idat[156]^idat[154]^idat[149]^idat[147]^idat[145]^idat[144]^idat[142]^idat[140]^idat[138]^idat[134]^idat[133]^idat[132]^idat[126]^idat[118]^idat[117]^idat[115]^idat[114]^idat[112]^idat[111]^idat[110]^idat[109]^idat[106]^idat[105]^idat[104]^idat[103]^idat[102]^idat[101]^idat[99]^idat[96]^idat[93]^idat[92]^idat[91]^idat[89]^idat[87]^idat[86]^idat[85]^idat[84]^idat[83]^idat[79]^idat[76]^idat[74]^idat[73]^idat[68]^idat[67]^idat[66]^idat[65]^idat[63]^idat[62]^idat[59]^idat[55]^idat[53]^idat[52]^idat[51]^idat[49]^idat[48]^idat[47]^idat[44]^idat[42]^idat[39]^idat[38]^idat[34]^idat[33]^idat[30]^idat[29]^idat[27]^idat[22]^idat[20]^idat[18]^idat[17]^idat[15]^idat[13]^idat[11]^idat[7]^idat[6]^idat[5]^icrc[5];

endmodule
