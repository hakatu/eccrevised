// megafunction wizard: %LPM_ADD_SUB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_ADD_SUB 

// ============================================================
// File Name: aladder.v
// Megafunction Name(s):
//          LPM_ADD_SUB
//
// Simulation Library Files(s):
//          lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
`define     RTL_SIMULATION
// synopsys translate_on
module aladder (
    cin,
    clock,
    dataa,
    datab,
    cout,
    result);

    input     cin;
    input     clock;
    input   [255:0]  dataa;
    input   [255:0]  datab;
    output    cout;
    output  [255:0]  result;

`ifndef RTL_SIMULATION

    wire  sub_wire0;
    wire [255:0] sub_wire1;
    wire  cout = sub_wire0;
    wire [255:0] result = sub_wire1[255:0];

    lpm_add_sub LPM_ADD_SUB_component (
                .cin (cin),
                .clock (clock),
                .dataa (dataa),
                .datab (datab),
                .cout (sub_wire0),
                .result (sub_wire1)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .clken (),
                .overflow ()
                // synopsys translate_on
                );
    defparam
        LPM_ADD_SUB_component.lpm_direction = "ADD",
        LPM_ADD_SUB_component.lpm_hint = "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=YES",
        LPM_ADD_SUB_component.lpm_pipeline = 2,
        LPM_ADD_SUB_component.lpm_representation = "UNSIGNED",
        LPM_ADD_SUB_component.lpm_type = "LPM_ADD_SUB",
        LPM_ADD_SUB_component.lpm_width = 256;

`else

reg [255:0] r;
reg         co;

always @(*)
    begin
    case(cin)
        1'b0: {co,r} = {1'b0,dataa} + {1'b0,datab};
        1'b1: {co,r} = {1'b0,dataa} - {1'b0,datab};
    endcase
    end

ffxkclkx #(2,256) u1 (clock, , r , result);
ffxkclkx #(2,1) u2 (clock, , co^cin , cout);

`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: CarryIn NUMERIC "1"
// Retrieval info: PRIVATE: CarryOut NUMERIC "1"
// Retrieval info: PRIVATE: ConstantA NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: Function NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "2"
// Retrieval info: PRIVATE: Latency NUMERIC "1"
// Retrieval info: PRIVATE: Overflow NUMERIC "0"
// Retrieval info: PRIVATE: RadixA NUMERIC "10"
// Retrieval info: PRIVATE: RadixB NUMERIC "10"
// Retrieval info: PRIVATE: Representation NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: ValidCtA NUMERIC "0"
// Retrieval info: PRIVATE: ValidCtB NUMERIC "0"
// Retrieval info: PRIVATE: WhichConstant NUMERIC "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: nBit NUMERIC "256"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: LPM_HINT STRING "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=YES"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "2"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_ADD_SUB"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "256"
// Retrieval info: USED_PORT: cin 0 0 0 0 INPUT NODEFVAL "cin"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: cout 0 0 0 0 OUTPUT NODEFVAL "cout"
// Retrieval info: USED_PORT: dataa 0 0 256 0 INPUT NODEFVAL "dataa[255..0]"
// Retrieval info: USED_PORT: datab 0 0 256 0 INPUT NODEFVAL "datab[255..0]"
// Retrieval info: USED_PORT: result 0 0 256 0 OUTPUT NODEFVAL "result[255..0]"
// Retrieval info: CONNECT: @cin 0 0 0 0 cin 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 256 0 dataa 0 0 256 0
// Retrieval info: CONNECT: @datab 0 0 256 0 datab 0 0 256 0
// Retrieval info: CONNECT: cout 0 0 0 0 @cout 0 0 0 0
// Retrieval info: CONNECT: result 0 0 256 0 @result 0 0 256 0
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL aladder_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
