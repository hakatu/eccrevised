////////////////////////////////////////////////////////////////////////////////
//
// Arrive Technologies
//
// Filename     : half_adder.v
// Description  : .
//
// Author       : hungnt@HW-NTHUNG
// Created On   : Tue Nov 06 11:40:02 2018
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module half_adder
    (
     a,
     b,
     sum,
     c
     );

////////////////////////////////////////////////////////////////////////////////
// Port declarations

input a;
input b;

output sum;
output c;

////////////////////////////////////////////////////////////////////////////////
// Output declarations

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations

////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation

assign sum = a ^ b;
assign c = a & b;

endmodule 
