////////////////////////////////////////////////////////////////////////////////
//
// Arrive Technologies
//
// Filename     : decodex.v
// Description  : Parameterized decoding from an number to a bitmap.
//
// Author       : lqcuong@HW-LQCUONG
// Created On   : Wed Jul 12 09:21:13 2006
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module decodex
    (
     in,
     out
     );

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations
parameter INWID = 6;
parameter OUTWID = 48;
parameter VALUE = 1'b1;

////////////////////////////////////////////////////////////////////////////////
// Port declarations
input [INWID-1:0] in;

output [OUTWID-1:0] out;

////////////////////////////////////////////////////////////////////////////////
// Output declarations


////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation

reg [OUTWID-1:0]    out;
always @(in)
begin
    out = {OUTWID{!VALUE}};
    out[in] = VALUE;
end

endmodule 
