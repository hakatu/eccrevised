module ATAND2
    (
     A,
     B,
     Y
     );
input A;
input B;
output Y;

wire   Y;
assign Y = A&B;

endmodule
//cao 