////////////////////////////////////////////////////////////////////////////////
//
// Arrive Technologies
//
// Filename     : ecc_enc16.v
// Description  : Encode 16 bits data using Hamming SEC code
//
// Author       : pmduc@HW-PMDUC
// Created On   : Mon Jun 05 14:45:19 2006
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module ecc_enc32
    (
     idat,
     odat    
     );
input   [31:0]   idat;
output  [37:0]   odat;
wire            p1,p2,p4,p8,p16,p32;
wire            d3,d5,d6,d7,d9,d10,d11,d12,d13,d14,d15,d17,d18,d19,d20,d21,
                d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d33,d34,d35,d36,d37,
                d38;

assign          {d38,d37,d36,d35,d34,d33,d31,d30,d29,d28,d27,d26,d25,d24,d23,d22,
                 d21,d20,d19,d18,d17,d15,d14,d13,d12,d11,d10,d9,d7,d6,d5,d3} = idat;

assign          p1 = d3 ^ d5 ^ d7 ^ d9 ^ d11 ^ d13 ^ d15 ^ d17 ^ d19 ^ d21 
                      ^ d23 ^ d25 ^ d27 ^ d29 ^ d31 ^ d33 ^ d35 ^ d37;

assign          p2 = d3 ^ d6 ^ d7 ^ d10 ^ d11 ^ d14 ^ d15 ^ d18 ^ d19 ^ d22 ^ 
                    d23 ^ d26 ^ d27 ^ d30 ^ d31 ^ d34 ^ d35 ^ d38;

assign          p4 = d5 ^ d6 ^ d7 ^ d12^ d13 ^ d14 ^ d15 ^ d20 ^ d21 ^ d22 ^ d23 ^
                    d28 ^ d29 ^ d30 ^ d31 ^ d36 ^ d37 ^ d38;

assign          p8 = d9 ^ d10^ d11^ d12^ d13 ^ d14 ^ d15 ^ d24 ^ d25 ^ d26 ^ d27 ^ 
                    d28 ^ d29 ^ d30 ^ d31;
assign          p16= d17 ^ d18 ^ d19 ^ d20 ^ d21 ^ d22 ^ d23 ^ d24 ^ d25 ^ d26 ^ d27 ^ d28 ^
                     d29 ^ d30 ^ d31;
assign          p32 = d33 ^ d34 ^ d35 ^ d36 ^ d37 ^ d38;


assign          odat = {d38,d37,d36,d35,d34,d33,p32,d31,d30,d29,d28,d27,d26,d25,d24,
                        d23,d22,d21,d20,d19,d18,d17,p16,d15,d14,d13,d12,d11,d10,d9,p8,d7,
                        d6,d5,p4,d3,p2,p1};
endmodule 

/*
-------------   p1  p2  p4  p8  p16  p32 p64
1   00001   p1                  
2   00010   p2                  
3   00011   d3  *   *           
4   00100   p4          *       
5   00101   d5  *       *   
6   00110   d6      *   *   
7   00111   d7  *   *   *       
8   01000   p8                  
9   01001   d9  *           *   
10  01010   d10     *       *   
11  01011   d11 *   *       *   
12  01100   d12         *   *   
13  01101   d13 *       *   *   
14  01110   d14     *   *   *   
15  01111   d15 *   *   *   *   
16  10000   p16                 
17  10001   d17 *               *
18  10010   d18     *           *
19  10011   d19 *   *           *
20  10100   d20         *       *
21  10101   d21 *       *       *
22  10110   d22     *   *       *
23  10111   d23 *   *   *       *
24  11000   d24             *   *
25  11001   d25 *           *   *
26  11010   d26     *       *   *
27  11011   d27 *   *       *   *
28  11100   d28         *   *   *
29  11101   d29 *       *   *   *
30  11110   d30     *   *   *   *
31  11111   d31 *   *   *   *   *
32 100000   p32                        
33 100001   d33 *                      *
34 100010   d34     *                  *
35 100011   d35 *   *                  *
36 100100   d36         *              *
37 100101   d37 *       *              *
38 100110   d38     *   *              *
39 100111   d39 *   *   *              *
40 101000   d40              *         *
41 101001   d41 *            *         *
42 101010   d42     *        *         *
43 101011   d43 *   *        *         *
44 101100   d44         *    *         *
45 101101   d45 *       *    *         *
46 101110   d46     *   *    *         *
47 101111   d47 *   *   *    *         *
48 110000   d48                  *     *
49 110001   d49 *                *     * 
50 110010   d50     *            *     *
51 110011   d51 *   *            *     *
52 110100   d52         *        *     * 
53 110101   d53 *       *        *     *
54 110110   d54     *   *        *     *
55 110111   d55 *   *   *        *     *
56 111000   d56              *   *     *
57 111001   d57 *            *   *     *
58 111010   d58     *        *   *     *
59 111011   d59 *   *        *   *     *
60 111100   d60         *    *   *     *
61 111101   d61 *       *    *   *     *
62 111110   d62     *   *    *   *     *
63 111111   d63 *   *   *    *   *     *
641000000   p64     
651000001   d65 *                           *
661000010   d66     *                       *
671000011   d67 *   *                       *
681000100   d68         *                   *
691000101   d69 *       *                   * 
701000110   d70     *   *                   *
711000111   d71 *   *   *                   *
*/  