module ippcrc_crc12_128b
    (
     ci,
     di,

     co
     );

////////////////////////////////////////////////////////////////////////////////
// Port declarations
input [11:0]   ci;
input [127:0]   di;

output [11:0]  co;

////////////////////////////////////////////////////////////////////////////////
// Output declarations
wire [11:0]    co;

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations

////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation
wire [11:0]     swdi;
assign          swdi =  {di[0],di[1],di[2],di[3],di[4],di[5],di[6],di[7],di[8],di[9],di[10],di[11]};

wire [11:0]     dx;
assign          dx   =  ci[11:0]^swdi[11:0];

assign          co[11]=dx[11]^dx[10]^dx[8]^dx[6]^dx[5]^dx[4]^
                di[13]^di[19]^di[20]^di[23]^di[26]^di[27]^di[32]^di[33]^di[34]^di[39]^di[40]^di[46]^di[47]^di[52]^di[53]^di[56]^di[58]^di[59]^di[62]^di[64]^di[65]^di[67]^di[68]^di[69]^di[70]^di[74]^di[76]^di[77]^di[78]^di[79]^di[80]^di[81]^di[84]^di[93]^di[94]^di[95]^di[98]^di[99]^di[102]^di[103]^di[104]^di[105]^di[106]^di[111]^di[112]^di[113]^di[114]^di[115]^di[116]^di[117]^di[120]^di[121]^di[122]^di[123]^di[124]^di[125]^di[126]^di[127];

assign          co[10]=dx[9]^dx[8]^dx[7]^dx[6]^dx[3]^
                di[13]^di[14]^di[19]^di[21]^di[23]^di[24]^di[26]^di[28]^di[32]^di[35]^di[39]^di[41]^di[46]^di[48]^di[52]^di[54]^di[56]^di[57]^di[58]^di[60]^di[62]^di[63]^di[64]^di[66]^di[67]^di[71]^di[74]^di[75]^di[76]^di[82]^di[84]^di[85]^di[93]^di[96]^di[98]^di[100]^di[102]^di[107]^di[111]^di[118]^di[120];

assign          co[9]=dx[11]^dx[8]^dx[7]^dx[6]^dx[5]^dx[2]^
                di[14]^di[15]^di[20]^di[22]^di[24]^di[25]^di[27]^di[29]^di[33]^di[36]^di[40]^di[42]^di[47]^di[49]^di[53]^di[55]^di[57]^di[58]^di[59]^di[61]^di[63]^di[64]^di[65]^di[67]^di[68]^di[72]^di[75]^di[76]^di[77]^di[83]^di[85]^di[86]^di[94]^di[97]^di[99]^di[101]^di[103]^di[108]^di[112]^di[119]^di[121];

assign          co[8]=dx[10]^dx[7]^dx[6]^dx[5]^dx[4]^dx[1]^
                di[15]^di[16]^di[21]^di[23]^di[25]^di[26]^di[28]^di[30]^di[34]^di[37]^di[41]^di[43]^di[48]^di[50]^di[54]^di[56]^di[58]^di[59]^di[60]^di[62]^di[64]^di[65]^di[66]^di[68]^di[69]^di[73]^di[76]^di[77]^di[78]^di[84]^di[86]^di[87]^di[95]^di[98]^di[100]^di[102]^di[104]^di[109]^di[113]^di[120]^di[122];

assign          co[7]=dx[11]^dx[9]^dx[6]^dx[5]^dx[4]^dx[3]^dx[0]^
                di[16]^di[17]^di[22]^di[24]^di[26]^di[27]^di[29]^di[31]^di[35]^di[38]^di[42]^di[44]^di[49]^di[51]^di[55]^di[57]^di[59]^di[60]^di[61]^di[63]^di[65]^di[66]^di[67]^di[69]^di[70]^di[74]^di[77]^di[78]^di[79]^di[85]^di[87]^di[88]^di[96]^di[99]^di[101]^di[103]^di[105]^di[110]^di[114]^di[121]^di[123];

assign          co[6]=dx[11]^dx[10]^dx[8]^dx[5]^dx[4]^dx[3]^dx[2]^
                di[12]^di[17]^di[18]^di[23]^di[25]^di[27]^di[28]^di[30]^di[32]^di[36]^di[39]^di[43]^di[45]^di[50]^di[52]^di[56]^di[58]^di[60]^di[61]^di[62]^di[64]^di[66]^di[67]^di[68]^di[70]^di[71]^di[75]^di[78]^di[79]^di[80]^di[86]^di[88]^di[89]^di[97]^di[100]^di[102]^di[104]^di[106]^di[111]^di[115]^di[122]^di[124];

assign          co[5]=dx[11]^dx[10]^dx[9]^dx[7]^dx[4]^dx[3]^dx[2]^dx[1]^
                di[13]^di[18]^di[19]^di[24]^di[26]^di[28]^di[29]^di[31]^di[33]^di[37]^di[40]^di[44]^di[46]^di[51]^di[53]^di[57]^di[59]^di[61]^di[62]^di[63]^di[65]^di[67]^di[68]^di[69]^di[71]^di[72]^di[76]^di[79]^di[80]^di[81]^di[87]^di[89]^di[90]^di[98]^di[101]^di[103]^di[105]^di[107]^di[112]^di[116]^di[123]^di[125];

assign          co[4]=dx[10]^dx[9]^dx[8]^dx[6]^dx[3]^dx[2]^dx[1]^dx[0]^
                di[14]^di[19]^di[20]^di[25]^di[27]^di[29]^di[30]^di[32]^di[34]^di[38]^di[41]^di[45]^di[47]^di[52]^di[54]^di[58]^di[60]^di[62]^di[63]^di[64]^di[66]^di[68]^di[69]^di[70]^di[72]^di[73]^di[77]^di[80]^di[81]^di[82]^di[88]^di[90]^di[91]^di[99]^di[102]^di[104]^di[106]^di[108]^di[113]^di[117]^di[124]^di[126];

assign          co[3]=dx[9]^dx[8]^dx[7]^dx[5]^dx[2]^dx[1]^dx[0]^
                di[12]^di[15]^di[20]^di[21]^di[26]^di[28]^di[30]^di[31]^di[33]^di[35]^di[39]^di[42]^di[46]^di[48]^di[53]^di[55]^di[59]^di[61]^di[63]^di[64]^di[65]^di[67]^di[69]^di[70]^di[71]^di[73]^di[74]^di[78]^di[81]^di[82]^di[83]^di[89]^di[91]^di[92]^di[100]^di[103]^di[105]^di[107]^di[109]^di[114]^di[118]^di[125]^di[127];

assign          co[2]=dx[10]^dx[7]^dx[5]^dx[1]^dx[0]^
                di[12]^di[16]^di[19]^di[20]^di[21]^di[22]^di[23]^di[26]^di[29]^di[31]^di[33]^di[36]^di[39]^di[43]^di[46]^di[49]^di[52]^di[53]^di[54]^di[58]^di[59]^di[60]^di[66]^di[67]^di[69]^di[71]^di[72]^di[75]^di[76]^di[77]^di[78]^di[80]^di[81]^di[82]^di[83]^di[90]^di[92]^di[94]^di[95]^di[98]^di[99]^di[101]^di[102]^di[103]^di[105]^di[108]^di[110]^di[111]^di[112]^di[113]^di[114]^di[116]^di[117]^di[119]^di[120]^di[121]^di[122]^di[123]^di[124]^di[125]^di[127];

assign          co[1]=dx[11]^dx[10]^dx[9]^dx[8]^dx[5]^dx[0]^
                di[12]^di[17]^di[19]^di[21]^di[22]^di[24]^di[26]^di[30]^di[33]^di[37]^di[39]^di[44]^di[46]^di[50]^di[52]^di[54]^di[55]^di[56]^di[58]^di[60]^di[61]^di[62]^di[64]^di[65]^di[69]^di[72]^di[73]^di[74]^di[80]^di[82]^di[83]^di[91]^di[94]^di[96]^di[98]^di[100]^di[105]^di[109]^di[116]^di[118]^di[127];

assign          co[0]=dx[11]^dx[9]^dx[7]^dx[6]^dx[5]^
                di[12]^di[18]^di[19]^di[22]^di[25]^di[26]^di[31]^di[32]^di[33]^di[38]^di[39]^di[45]^di[46]^di[51]^di[52]^di[55]^di[57]^di[58]^di[61]^di[63]^di[64]^di[66]^di[67]^di[68]^di[69]^di[73]^di[75]^di[76]^di[77]^di[78]^di[79]^di[80]^di[83]^di[92]^di[93]^di[94]^di[97]^di[98]^di[101]^di[102]^di[103]^di[104]^di[105]^di[110]^di[111]^di[112]^di[113]^di[114]^di[115]^di[116]^di[119]^di[120]^di[121]^di[122]^di[123]^di[124]^di[125]^di[126]^di[127];


endmodule