// megafunction wizard: %ALTDDIO_OUT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altddio_out 

// ============================================================
// File Name: alt_ddr_output.v
// Megafunction Name(s):
//          altddio_out
//
// Simulation Library Files(s):
//          altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Build 151 09/26/2007 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
//`timescale 1 ps / 1 ps
// synopsys translate_on
module alt_ddr_output (
    datain_h,
    datain_l,
    outclock,
    dataout);

parameter   PAD_WIDTH = 8;

    input   [PAD_WIDTH-1:0]  datain_h;
    input   [PAD_WIDTH-1:0]  datain_l;
    input     outclock;
    output  [PAD_WIDTH-1:0]  dataout;

wire [PAD_WIDTH-1:0]         dataout;
assign                       dataout = outclock ? datain_h : datain_l;

endmodule
